*----------------------------------------------------------------------
* res_mp.cir
*
* SPICE Netlist: Resistor with multiple parameters
*
* Copyright(C) 2014 MetaMorph Inc.
* http://metamorphsoftware.com/
*
*
*----------------------------------------------------------------------
*----------------------------------------------------------------------
* 
* 
* 
*        (1)
*         o-----------.
*                     |
*                     | L1
*                     C|
*                     C|
*                     C|
*                     |
*                     | (11)
*                     |
*                     |
*                     | R1
*                    .-.
*                    | |
*                    | |
*                    '-'
*                     |
*        (2)          |
*         o-----------'
* 
* 
*   
*----------------------------------------------------------------------
.SUBCKT RES_MP 1 2 RVAL=1.0k LVAL=800pH
L1  1 11 LVAL
R1 11  2 RVAL
.ENDS RES_MP


