*----------------------------------------------------------------------
* res_0603_330R.cir
*
* SPICE Netlist: Resistor chip, 0603 package, 330 Ohms
*
* Copyright(C) 2014 MetaMorph Inc.
* http://metamorphsoftware.com/
*
*
*----------------------------------------------------------------------
*----------------------------------------------------------------------
* 
* 
* 
*        (1)
*         o-----------.
*                     |
*                     |
*                     | R1
*                    .-.
*                    | |
*                    | |
*                    '-'
*                     |
*        (2)          |
*         o-----------'
* 
* 
*   
*----------------------------------------------------------------------
.MODEL RES_0603_330 R RES=1.0k


